module counter_top (
    input logic sysclk,
    output logic [3:0] led
);
  logic clksel, clkpulse, clkout, rst, load, up_down, enable;
  logic [3:0] d_in, count;

  // Select the clock
  assign clkout = (clksel) ? sysclk : clkpulse;
  assign led = count;

  // Instantiate DUT
  updown_counter dut0 (
      .clk    (clkout),
      .rst  (rst),
      //.load   (load),     // Load enable
      .up_down(up_down),  // Direction control (1 = up, 0 = down)
      .enable (enable),   // Counter enable
      //.d_in   (d_in),     // Input data for loading
      .count  (count)     // Counter output
  );
//  updown_counter dut0 (
//      .clk    (clkout),
//      .rst_n  (1'b1),
//      .load   (1'b1),     // Load enable
//      .up_down(1'b1),  // Direction control (1 = up, 0 = down)
//      .enable (1'b1),   // Counter enable
//      .d_in   (4'b0000),     // Input data for loading
//      .count  (count)     // Counter output
//  );

  // VIO for control signals
    vio_0 vio0 (
      .clk(sysclk),  // Use actual clock
      .probe_out0(clksel),
      .probe_out1(clkpulse),
      .probe_out2(rst),
      //.probe_out3(load),
      .probe_out3(up_down),
      .probe_out4(enable),
     // .probe_out6(d_in),
      .probe_in0(count)
  );

    // ILA to monitor counter output in free running mode
    // Also takes in the enable so triggering can be demonstrated
    ila_0 ila0 (
        .clk(sysclk), // Actual system clock
        .probe0(enable),
        .probe1(count)
    );

endmodule
